module top_module(output reg one);
	assign one = 1'b1
endmodule